module ins_mem(ins_out,add,rst);
input [31:0]add;
input rst;
output reg [31:0]ins_out;
reg [31:0]mem[255:0];

always@(*)
begin
    if(rst==1)
    begin
        // add
        mem[0] = 32'b00000000010111000000110010110011;
        // sub
        mem[1] = 32'b01100000001100110000000101011011;
        // lw
        
        mem[2] = 32'b0000000000000000010000101100000;
        mem[3] = 32'b00000000000101001000010010010011;
        mem[4] = 32'b00000000010111000000110010110011;
        mem[5] = 32'b00100100000100010000000000001011;
        mem[6] = 32'b00000000000100010000000100000011;
        mem[7] =32'b01000000000100010000000100000011;
        mem[8] =  32'b00000000000100010000000111100111;
        mem[9] =  32'b00000000001000010000100010000011;
        mem[10] =  32'b00000000000000010000000000001011;
        mem[11] =  32'b00000000000000010000000000001011;
        mem[12] = 32'b00000000000000010000000000001011;
        mem[13] =  32'b01000000000100010000000000100011;
        mem[14] =  32'b00000000000100010000000000100011;
        mem[15] =   32'b00100100001100010000000000010100;
        mem[16] =  32'b00000000001100010000000100000011;
        mem[17] =  32'b01000000001100010000000100000011;
        mem[18] =  32'b00000000001100010000000111100111;
        mem[19] =  32'b00000000001100010000000111000111;
        mem[20] =  32'b00000000000000100000000000010100;
        mem[21] =  32'b00000000000000100000000000010100;
        mem[22] =  32'b00000000000000100000000000010100;
        mem[23] =  32'b01000000001100010000000001010011;
        mem[24] =  32'b00000000001100010000000001010011;
        mem[25] =   32'b00100100010100010000000000011110;
        mem[26] =  32'b0000000001010001000000010000011;
        mem[27] =  32'b0100000001010001000000010000011;
        mem[28] =   32'b00000000010100010000000111100111;
        mem[29] =   32'b00000000010100010000000111000111;
        mem[30] =   32'b00000000000000011000000000011110;
        mem[31] =   32'b00000000000000011000000000011110;
        mem[32] =   32'b00000000000000011000000000011110;
        mem[33] =   32'b01000000010100010000000001111011;
        mem[34] =   32'b00000000010100010000000001111011;
        mem[35] =  32'b00100100100001110000000000101000;
        mem[36] =  32'b00000000001001110000100100000011;
    end
    ins_out = mem[add];
end
endmodule